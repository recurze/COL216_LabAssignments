package mytypes is
	type state is (fetch,rdAB,arith,wrRF,addr,wrM,rdM,M2RF,brn,nope);
end package;
package body mytypes is
end mytypes;
